clkDIV